entity or_gate is
  port (
    a, b : in bit;
    q : out bit
  );  
end entity;

architecture structural of or_gate is
begin
end structural;

--

entity or_gate_tb is
end entity;

architecture behavior of or_gate_tb is
begin

end architecture;
